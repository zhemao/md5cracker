module md5cracker (
    input clock_50,
    output [3:0] leds
);

endmodule